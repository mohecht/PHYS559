* Qubit Energy Tuner

.model jj1 jj(level=1)

.control
run
plot .
save .
.endc



B1 1 15 100 jj1 ics=160uA 
B2 5 17 100 jj1 ics=160uA 
B3 8 19 100 jj1 ics=160uA
B4 12 21 100 jj1 ics=160uA
K1 L4 LN4 .08
K2 L3 LN3 .08
K3 L2 LN2 .8
K4 L1 LN1 .8
L1 1 0 10nH
L2 0 5 10nH
L3 8 0 10nH
L4 0 12 10nH
L11 15 4 0.05pH
L12 16 4 0.955pH
L13 4 0 0.096pH
L21 17 7 0.05pH
L22 18 7 0.955pH
L23 7 0 0.096pH
L31 19 11 0.05pH
L32 20 11 0.955pH
L33 11 0 0.096pH
L41 21 14 0.05pH
L42 22 14 0.955pH
L43 14 0 0.096pH
LN0 10 0 1nH
LN1 2 3 10nH
LN2 3 6 10nH
LN3 6 9 10nH
LN4 9 13 10nH
LN5 13 10 2nH
R1 1 16 0.766
R2 5 18 0.766
R3 8 20 0.766
R4 12 22 0.766
VA 1 0 gpulse(0 0 20ps 1ps)+ gpulse(0 0 100ps 1ps)+gpulse(0 0 120ps 1ps)+gpulse(0 0 300ps 1ps)+gpulse(0 0 380ps 1ps)+gpulse(0 0 400ps 1ps)
VB 5 0 gpulse(0 0 40ps 1ps)+gpulse(0 0 180ps 1ps)+gpulse(0 0 200ps 1ps) +gpulse(0 0 360ps 1ps)+gpulse(0 0 420ps 1ps)+gpulse(0 0 440ps 1ps)
VC 8 0 gpulse(0 0 60ps 1ps)+gpulse(0 0 140ps 1ps)+gpulse(0 0 220ps 1ps)+gpulse(0 0 240ps 1ps)+gpulse(0 0 320ps  1ps)
VD 12 0 gpulse(0 0 80ps 1ps)+gpulse(0 0 160ps 1ps)+gpulse(0 0 260ps 1ps)+gpulse(0 0 280ps 1ps)+gpulse(0 0 340ps 1ps)
VP0 2 0


.tran .005p 460ps uic

.plot tran @VP0[c] v(1) v(5) v(8) v(12) 


.save tran
.save v(12) 
.save v(8) 
.save @VP0[c]
.save v(5)
.save v(1)

** C:\Users\malid\qet.cir

