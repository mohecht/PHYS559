.model jj0 jj(rtype = 2 icrit=225uA cap=450.0000fF)
.model jj1 jj(rtype = 2 icrit=250uA cap=600.0000fF)
.model jj2 jj(rtype = 2 icrit=160uA cap=600.0000fF)



IA 2 0 pulse(0uA 300uA 2ns 0.01ns 0.01ns 1ns)
IB 14 0 pulse(0uA 300uA 4ns 0.01ns 0.01ns 1ns)
IC 25 0 pulse(0uA 300uA 6ns 0.01ns 0.01ns 1ns)
ID 37 0 pulse(0uA 300uA 10ns 0.01ns 0.01ns 1ns)
BJ1 8 54 0 jj2 
BJ2 19 65 0 jj2 
BJ3 30 76 0 jj2 
BJ4 42 87 0 jj2 
BJJ1A 5 49 0 jj0 
BJJ1B 16 60 0 jj0 
BJJ1C 27 71 0 jj0 
BJJ1D 39 82 0 jj0 
BJJ2A 6 50 0 jj0
BJJ2B 17 61 0 jj0
BJJ2C 28 72 0 jj0 
BJJ2D 40 83 0 jj0 
BJJ3A 7 52 0 jj1 
BJJ3B 18 63 1000 jj1 
BJJ3C 29 74 0 jj1 
BJJ3D 41 85 0 jj1 
K1 L4 LN4 0.08
K2 L1 LN1 0.8
K3 L2 LN2 0.8
K4 L3 LN3 0.08
K5 L1 L2 0.7023
K6 L3 L4 0.7023
L1 8 0 10nH
L2 19 0 10nH
L3 30 0 10nH
L4 42 0 10nH
L11 54 12 0.05pH
L12 55 12 0.955pH
L13 12 0 0.096pH
L21 65 23 0.05pH
L22 66 23 0.955pH
L23 23 0 0.096pH
L31 76 35 0.05pH
L32 77 35 0.955pH
L33 35 0 0.096pH
L41 87 46 0.05pH
L42 88 46 0.955pH
L43 46 0 0.096pH
LJ11A 49 4 0.058pH
LJ11B 60 15 0.058pH
LJ11C 71 26 0.058pH
LJ11D 82 38 0.058pH
LJ12A 56 4 0.945pH
LJ12B 67 15 0.945pH
LJ12C 78 26 0.945pH
LJ12D 89 38 0.945pH
LJ13A 3 4 0.355pH
LJ13C 70 26 0.355pH
LJ13D 81 38 0.355pH
LJ21A 50 10 0.05pH
LJ21B 61 21 0.05pH
LJ21C 72 33 0.05pH
LJ21D 83 44 0.05pH
LJ22A 51 10 0.955pH
LJ22B 62 21 0.955pH
LJ22C 73 33 0.955pH
LJ22D 84 44 0.955pH
LJ23A 10 0 0.096pH
LJ23B 21 0 0.096pH
LJ23C 33 0 0.096pH
LJ23D 44 0 0.096pH
LJ31A 52 11 0.028pH
LJ31B 63 22 0.028pH
LJ31C 74 34 0.028pH
LJ31D 85 45 0.028pH
LJ32A 53 11 0.961pH
LJ32B 64 22 0.961pH
LJ32C 75 34 0.961pH
LJ32D 86 45 0.961pH
LJ33A 11 0 0.103pH
LJ33B 22 0 0.103pH
LJ33C 34 0 0.103pH
LJ33D 45 0 0.103pH
LN0 32 0 1nH
LN1 0 9 10nH
LN2 9 20 10nH
LN3 20 31 10nH
LN4 31 43 10nH
LN5 43 32 2nH
LQ1A 2 3 1.071pH
LQ1B 14 59 1.071pH
LQ1C 25 70 1.071pH
LQ1D 37 81 1.071pH
LQ2A 3 0 3.927pH
LQ2B 59 0 3.927pH
LQ2C 70 0 3.927pH
LQ2D 81 0 3.927pH
LQ3A 5 6 0.913pH
LQ3B 16 17 0.913pH
LQ3C 27 28 0.913pH
LQ3D 39 40 0.913pH
LQ4A 6 7 4.399pH
LQ4B 17 18 4.399pH
LQ4C 28 29 4.399pH
LQ4D 40 41 4.399pH
LQ5A 7 8 1.09pH
LQ5B 18 19 1.09pH
LQ5C 29 30 1.090pH
LQ5D 41 42 1.09pH
LV1A 47 5 16.8pH
LV1B 57 16 16.8pH
LV1C 68 27 16.8pH
LV1D 79 39 16.8pH
LV2A 48 7 15.5pH
LV2B 58 18 15.5pH
LV2C 69 29 15.5pH
LV2D 80 41 15.5pH
R1 8 55 0.766
R2 19 66 0.766
R3 30 77 0.766
R4 42 88 0.766
RJ1A 5 56 0.766
RJ1B 16 67 0.766
RJ1C 27 78 0.766
RJ1D 39 89 0.766
RJ2A 6 51 0.766
RJ2B 17 62 0.766
RJ2C 28 73 0.766
RJ2D 40 84 0.766
RJ3B 18 64 0.688
RJ3C 29 75 0.688
RJ3D 41 86 0.688
RV1A 1 47 9.09
RV1B 13 57 9.09
RV1C 24 68 9.09
RV1D 36 79 9.09
RV2A 1 48 14.29
RV2B 13 58 14.29
RV2C 24 69 14.29
RV2D 36 80 14.29
VQA 1 0 2.5mV
VQB 13 0 2.5mV
VQC 24 0 2.5mV
VQD 36 0 2.5mV
I_LN1 LN1 0 DC 0
* voltage nodes
VA 7 0 0V
VB 18 0 0V
VC 29 0 0V
VD 41 0 0V


.tran 0.05n 15n uic

.save @IA[c]
.save @IB[c]
.save @IC[c]
.save @ID[c]
.save V(7)
.save V(18)
.save V(29)
.save V(41)
.save I_LN1
